library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
entity InstructionMemory is
    Port ( rst : in  STD_LOGIC;
           address : in  STD_LOGIC_VECTOR (31 downto 0);
           imout : out  STD_LOGIC_VECTOR (31 downto 0):=(others=>'0'));
end InstructionMemory;
architecture Behavioral of InstructionMemory is
type rom_type is array (63 downto 0) of STD_LOGIC_VECTOR (31 downto 0);                 
	 signal ROM : rom_type:= (
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "10011000001000000100000000000010","10010110001110000100000000000010",
									  "10010100001010000100000000000010","10010010000110000100000000000010",
									  "10010000000000000100000000000010","10000100000100000011111111111001",
									  "10000010000100000010000000001000","00000001000000000000000000000000");
	signal rdata : std_logic_vector (31 downto 0);
begin
	rdata <= ROM(conv_integer(address));
	process (rst,address)
	begin
		  if (rst = '1') then
				imout <= ROM(conv_integer("00000000000000000000000000000000"));
		  else
				imout <= rdata;
		  end if;
	end process;
end Behavioral;